Dynamic Array in SystemVerilog :
 -As name dynamic suggests, an array whose size can be changed during run time simulation.
 -The size of an array can be specified during run-time by using new[ ]. 
 -Note: By default, the size of a dynamic array is 0 unless a new[ ] is used.
 -Hence ,Dynamic array is a concept ,where the space does not exist,untill the array is explicetely created during run time.
 -Dynamic array is an unpacked array whose sizes can be changed during run time.
 -The methods used in dynamic array are : new[] , size(), delete()


