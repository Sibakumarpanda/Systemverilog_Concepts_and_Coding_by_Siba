2_difference_between_@(event)_and_wait_(event.triggered)_with_example
