Array Locator methods :
