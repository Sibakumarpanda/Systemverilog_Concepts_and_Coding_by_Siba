Array reduction methods Overview :
  -The array reduction methods are used to reduce the array to a single value with the optional use of the ‘with’ clause.
  -The reduction methods can be applied on any unpacked array. 
  -For a ‘with’ clause, boolean or arithmetic reduction operation must be specified.
  -Note: If the ‘with’ clause is specified, the above reduction methods return value based on evaluating the expression for each array element.

Methods                                                     Description

and                                                         Returns bitwise AND (&) of all elements of the array.

or                                                          Returns bitwise OR (|) of all elements of the array.

xor                                                         Returns bitwise XOR (^) of all elements of the array.

sum                                                         Returns the sum of all elements of the array.

product                                                     Returns product of all elements of the array.

/**********************************************/
    Array Reduction Method Example1
/**********************************************/    
