SystemVerilog Queue Overview:
