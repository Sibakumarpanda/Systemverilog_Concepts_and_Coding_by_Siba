Array ordering methods in SV
  -The ordering methods are used to reorder the single-dimensional arrays or queues.

Methods                                                      Description

shuffle                                                      Randomizes the order of the elements in an array

sort                                                         Sorts the unpacked array in ascending order

rsort                                                        Sorts the unpacked array in descending order

reverse                                                      Reverses all the elements of a packed or unpacked array.
