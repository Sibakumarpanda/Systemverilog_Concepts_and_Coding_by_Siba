SystemVerilog Arrays :
 -An array is a group of variables having the same data type. It can be accessed using an index value. 
 -An index is a memory address and the array value is stored at that address.
Types of an array:
  1. Fixed-size array in SystemVerilog
  2. Single dimensional array
  3. Multidimensional array
     a. Two-dimensional array.
     b. Three-dimensional array
 4.  Packed and Unpacked array in SystemVerilog
 5.  Dynamic array in SystemVerilog
 6.  Associative array in SystemVerilog
